module SPIMaster(
    input i_clk,
    input i_reset
);

always @(posedge i_clk or posedge i_reset)
begin
end

endmodule
